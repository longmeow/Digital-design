`include "alu.v"

module alu_tb ();
    reg [31:0] a, b; //32-bit input
    reg [2:0] alu_sel; // 3-bit selection
    wire [31:0] alu_out; // 32-bit output
    wire carry_out;

    
endmodule